200000 2356 700 28 28 192 4 1
1 1 0 1 1 64
2 1 0 1 1 96
2 2 0 3 3 128
3 1 0 1 1 16
3 2 0 5 5 32
4 1 1 3 3 32
4 2 0 1 1 32